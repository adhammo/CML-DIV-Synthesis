.include dff_params.cir
.include dff.cir

.lib _PDK_ROOT/libs.tech/combined/sky130.lib.spice _CORNER

Xdff VDD VSS ip in op on ckp ckn dff winp={winp} wclk={wclk} wlat={wlat}
                                    +nfinp={nfinp} nfclk={nfclk} nflat={nflat}
                                    +vsw={vsw} iss={iss}

C1 op VSS {cload} m=1
C2 on VSS {cload} m=1

Xbalun1 indiff incm ip in balun
Xbalun2 clkdiff clkcm ckp ckn balun

vvdd VDD 0 1.8
vvss VSS 0 0
vinput indiff 0 dc {vsw_in} PULSE({-vsw_in} {vsw_in} 0 5p 5p 400p 800p)
vclk clkdiff 0 dc {vsw_clk} PULSE({-vsw_clk} {vsw_clk} 30p 5p 5p 400p 800p)
V1 incm 0 {1.8-vsw_in/2}
V2 clkcm 0 {1.8-cm_clk-vsw_clk/2}

.IC V(op)={1.8-vsw}
.IC V(on)={1.8}

.control

save all

set filetype = ascii
set hcopydevtype = svg
set format = cross

set appendwrite
echo "prop_delay" > outputs.csv

tran 1p 400p
let x = v(ckp)-v(ckn)
let y = v(op)-v(on)
meas tran tdiff TRIG x VAL=0 RISE=1 TARG y VAL=0 RISE=1

echo "$&tdiff" >> outputs.csv

.endc

.subckt balun d c p n
E1 net4 c d 0 0.5
V1 p net4 0
F1 d 0 V1 -0.5
R1 d 0 1T m=1
E2 net2 n d 0 0.5
V2 c net3 0
F2 d 0 V2 -0.5
R2 net3 net2 1u m=1
.ends

.end
