.param and_win1=$and_win1
.param and_win2=$and_win2
.param and_nfin1=$and_nfin1
.param and_nfin2=$and_nfin2
.param and_vsw=$and_vsw
.param and_iss=$and_iss
.param dff1_latch1_winp=$dff1_latch1_winp
.param dff1_latch1_wclk=$dff1_latch1_wclk
.param dff1_latch1_wlat=$dff1_latch1_wlat
.param dff1_latch1_nfinp=$dff1_latch1_nfinp
.param dff1_latch1_nfclk=$dff1_latch1_nfclk
.param dff1_latch1_nflat=$dff1_latch1_nflat
.param dff1_latch1_vsw=$dff1_latch1_vsw
.param dff1_latch1_iss=$dff1_latch1_iss
.param dff1_latch2_winp=$dff1_latch2_winp
.param dff1_latch2_wclk=$dff1_latch2_wclk
.param dff1_latch2_wlat=$dff1_latch2_wlat
.param dff1_latch2_nfinp=$dff1_latch2_nfinp
.param dff1_latch2_nfclk=$dff1_latch2_nfclk
.param dff1_latch2_nflat=$dff1_latch2_nflat
.param dff1_latch2_vsw=$dff1_latch2_vsw
.param dff1_latch2_iss=$dff1_latch2_iss
.param or_win1=$or_win1
.param or_win2=$or_win2
.param or_nfin1=$or_nfin1
.param or_nfin2=$or_nfin2
.param or_vsw=$or_vsw
.param or_iss=$or_iss
.param dff2_latch1_winp=$dff2_latch1_winp
.param dff2_latch1_wclk=$dff2_latch1_wclk
.param dff2_latch1_wlat=$dff2_latch1_wlat
.param dff2_latch1_nfinp=$dff2_latch1_nfinp
.param dff2_latch1_nfclk=$dff2_latch1_nfclk
.param dff2_latch1_nflat=$dff2_latch1_nflat
.param dff2_latch1_vsw=$dff2_latch1_vsw
.param dff2_latch1_iss=$dff2_latch1_iss
.param dff2_latch2_winp=$dff2_latch2_winp
.param dff2_latch2_wclk=$dff2_latch2_wclk
.param dff2_latch2_wlat=$dff2_latch2_wlat
.param dff2_latch2_nfinp=$dff2_latch2_nfinp
.param dff2_latch2_nfclk=$dff2_latch2_nfclk
.param dff2_latch2_nflat=$dff2_latch2_nflat
.param dff2_latch2_vsw=$dff2_latch2_vsw
.param dff2_latch2_iss=$dff2_latch2_iss
.param sf_w=$sf_w
.param sf_nf=$sf_nf
.param sf_iss=$sf_iss
.param vsw_clk=$vsw_clk
.param vsw_mc=$vsw_mc
.param cm_clk=$cm_clk
.param cwire=$cwire
.param cload=$cload