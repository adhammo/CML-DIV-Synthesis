.subckt divider VSS VDD op on ckp ckn latch1_winp=10 latch1_wclk=10 latch1_wlat=10 latch1_nfinp=5 latch1_nfclk=5 latch1_nflat=5 latch1_vsw=0.3 latch1_iss=1m latch2_winp=10 latch2_wclk=10 latch2_wlat=10 latch2_nfinp=5 latch2_nfclk=5 latch2_nflat=5 latch2_vsw=0.3 latch2_iss=1m sf_w=10 sf_nf=5 sf_iss=1m cwire=10f vdd=1.8
*.iopin VSS
*.iopin VDD
*.opin op
*.opin on
*.ipin ckp
*.ipin ckn

XM2 mn oin net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W={latch1_winp} nf={latch1_nfinp} ad='int(({latch1_nfinp} + 1)/2) * {latch1_winp} / {latch1_nfinp} * 0.29'
+ as='int(({latch1_nfinp} + 2)/2) * {latch1_winp} / {latch1_nfinp} * 0.29' pd='2*int(({latch1_nfinp} + 1)/2) * ({latch1_winp} / {latch1_nfinp} + 0.29)'
+ ps='2*int(({latch1_nfinp} + 2)/2) * ({latch1_winp} / {latch1_nfinp} + 0.29)' nrd='0.29 / {latch1_winp} ' nrs='0.29 / {latch1_winp} '
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 mp oip net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W={latch1_winp} nf={latch1_nfinp} ad='int(({latch1_nfinp} + 1)/2) * {latch1_winp} / {latch1_nfinp} * 0.29'
+ as='int(({latch1_nfinp} + 2)/2) * {latch1_winp} / {latch1_nfinp} * 0.29' pd='2*int(({latch1_nfinp} + 1)/2) * ({latch1_winp} / {latch1_nfinp} + 0.29)'
+ ps='2*int(({latch1_nfinp} + 2)/2) * ({latch1_winp} / {latch1_nfinp} + 0.29)' nrd='0.29 / {latch1_winp} ' nrs='0.29 / {latch1_winp} '
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 ckn net2 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W={latch1_wclk} nf={latch1_nfclk} ad='int(({latch1_nfclk} + 1)/2) * {latch1_wclk} / {latch1_nfclk} * 0.29'
+ as='int(({latch1_nfclk} + 2)/2) * {latch1_wclk} / {latch1_nfclk} * 0.29' pd='2*int(({latch1_nfclk} + 1)/2) * ({latch1_wclk} / {latch1_nfclk} + 0.29)'
+ ps='2*int(({latch1_nfclk} + 2)/2) * ({latch1_wclk} / {latch1_nfclk} + 0.29)' nrd='0.29 / {latch1_wclk} ' nrs='0.29 / {latch1_wclk} '
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net3 ckp net2 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W={latch1_wclk} nf={latch1_nfclk} ad='int(({latch1_nfclk} + 1)/2) * {latch1_wclk} / {latch1_nfclk} * 0.29'
+ as='int(({latch1_nfclk} + 2)/2) * {latch1_wclk} / {latch1_nfclk} * 0.29' pd='2*int(({latch1_nfclk} + 1)/2) * ({latch1_wclk} / {latch1_nfclk} + 0.29)'
+ ps='2*int(({latch1_nfclk} + 2)/2) * ({latch1_wclk} / {latch1_nfclk} + 0.29)' nrd='0.29 / {latch1_wclk} ' nrs='0.29 / {latch1_wclk} '
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 mn mp net3 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W={latch1_wlat} nf={latch1_nflat} ad='int(({latch1_nflat} + 1)/2) * {latch1_wlat} / {latch1_nflat} * 0.29'
+ as='int(({latch1_nflat} + 2)/2) * {latch1_wlat} / {latch1_nflat} * 0.29' pd='2*int(({latch1_nflat} + 1)/2) * ({latch1_wlat} / {latch1_nflat} + 0.29)'
+ ps='2*int(({latch1_nflat} + 2)/2) * ({latch1_wlat} / {latch1_nflat} + 0.29)' nrd='0.29 / {latch1_wlat} ' nrs='0.29 / {latch1_wlat} '
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 mp mn net3 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W={latch1_wlat} nf={latch1_nflat} ad='int(({latch1_nflat} + 1)/2) * {latch1_wlat} / {latch1_nflat} * 0.29'
+ as='int(({latch1_nflat} + 2)/2) * {latch1_wlat} / {latch1_nflat} * 0.29' pd='2*int(({latch1_nflat} + 1)/2) * ({latch1_wlat} / {latch1_nflat} + 0.29)'
+ ps='2*int(({latch1_nflat} + 2)/2) * ({latch1_wlat} / {latch1_nflat} + 0.29)' nrd='0.29 / {latch1_wlat} ' nrs='0.29 / {latch1_wlat} '
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 oin mp net5 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W={latch2_winp} nf={latch2_nfinp} ad='int(({latch2_nfinp} + 1)/2) * {latch2_winp} / {latch2_nfinp} * 0.29'
+ as='int(({latch2_nfinp} + 2)/2) * {latch2_winp} / {latch2_nfinp} * 0.29' pd='2*int(({latch2_nfinp} + 1)/2) * ({latch2_winp} / {latch2_nfinp} + 0.29)'
+ ps='2*int(({latch2_nfinp} + 2)/2) * ({latch2_winp} / {latch2_nfinp} + 0.29)' nrd='0.29 / {latch2_winp} ' nrs='0.29 / {latch2_winp} '
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 oip mn net5 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W={latch2_winp} nf={latch2_nfinp} ad='int(({latch2_nfinp} + 1)/2) * {latch2_winp} / {latch2_nfinp} * 0.29'
+ as='int(({latch2_nfinp} + 2)/2) * {latch2_winp} / {latch2_nfinp} * 0.29' pd='2*int(({latch2_nfinp} + 1)/2) * ({latch2_winp} / {latch2_nfinp} + 0.29)'
+ ps='2*int(({latch2_nfinp} + 2)/2) * ({latch2_winp} / {latch2_nfinp} + 0.29)' nrd='0.29 / {latch2_winp} ' nrs='0.29 / {latch2_winp} '
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 net5 ckp net6 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W={latch2_wclk} nf={latch2_nfclk} ad='int(({latch2_nfclk} + 1)/2) * {latch2_wclk} / {latch2_nfclk} * 0.29'
+ as='int(({latch2_nfclk} + 2)/2) * {latch2_wclk} / {latch2_nfclk} * 0.29' pd='2*int(({latch2_nfclk} + 1)/2) * ({latch2_wclk} / {latch2_nfclk} + 0.29)'
+ ps='2*int(({latch2_nfclk} + 2)/2) * ({latch2_wclk} / {latch2_nfclk} + 0.29)' nrd='0.29 / {latch2_wclk} ' nrs='0.29 / {latch2_wclk} '
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 net7 ckn net6 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W={latch2_wclk} nf={latch2_nfclk} ad='int(({latch2_nfclk} + 1)/2) * {latch2_wclk} / {latch2_nfclk} * 0.29'
+ as='int(({latch2_nfclk} + 2)/2) * {latch2_wclk} / {latch2_nfclk} * 0.29' pd='2*int(({latch2_nfclk} + 1)/2) * ({latch2_wclk} / {latch2_nfclk} + 0.29)'
+ ps='2*int(({latch2_nfclk} + 2)/2) * ({latch2_wclk} / {latch2_nfclk} + 0.29)' nrd='0.29 / {latch2_wclk} ' nrs='0.29 / {latch2_wclk} '
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 oin oip net7 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W={latch2_wlat} nf={latch2_nflat} ad='int(({latch2_nflat} + 1)/2) * {latch2_wlat} / {latch2_nflat} * 0.29'
+ as='int(({latch2_nflat} + 2)/2) * {latch2_wlat} / {latch2_nflat} * 0.29' pd='2*int(({latch2_nflat} + 1)/2) * ({latch2_wlat} / {latch2_nflat} + 0.29)'
+ ps='2*int(({latch2_nflat} + 2)/2) * ({latch2_wlat} / {latch2_nflat} + 0.29)' nrd='0.29 / {latch2_wlat} ' nrs='0.29 / {latch2_wlat} '
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 oip oin net7 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W={latch2_wlat} nf={latch2_nflat} ad='int(({latch2_nflat} + 1)/2) * {latch2_wlat} / {latch2_nflat} * 0.29'
+ as='int(({latch2_nflat} + 2)/2) * {latch2_wlat} / {latch2_nflat} * 0.29' pd='2*int(({latch2_nflat} + 1)/2) * ({latch2_wlat} / {latch2_nflat} + 0.29)'
+ ps='2*int(({latch2_nflat} + 2)/2) * ({latch2_wlat} / {latch2_nflat} + 0.29)' nrd='0.29 / {latch2_wlat} ' nrs='0.29 / {latch2_wlat} '
+ sa=0 sb=0 sd=0 mult=1 m=1
XM13 VDD oip op VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W={sf_w} nf={sf_nf} ad='int(({sf_nf} + 1)/2) * {sf_w} / {sf_nf} * 0.29' as='int(({sf_nf} + 2)/2) * {sf_w} / {sf_nf} * 0.29'
+ pd='2*int(({sf_nf} + 1)/2) * ({sf_w} / {sf_nf} + 0.29)' ps='2*int(({sf_nf} + 2)/2) * ({sf_w} / {sf_nf} + 0.29)' nrd='0.29 / {sf_w} '
+ nrs='0.29 / {sf_w} ' sa=0 sb=0 sd=0 mult=1 m=1
XM14 VDD oin on VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W={sf_w} nf={sf_nf} ad='int(({sf_nf} + 1)/2) * {sf_w} / {sf_nf} * 0.29' as='int(({sf_nf} + 2)/2) * {sf_w} / {sf_nf} * 0.29'
+ pd='2*int(({sf_nf} + 1)/2) * ({sf_w} / {sf_nf} + 0.29)' ps='2*int(({sf_nf} + 2)/2) * ({sf_w} / {sf_nf} + 0.29)' nrd='0.29 / {sf_w} '
+ nrs='0.29 / {sf_w} ' sa=0 sb=0 sd=0 mult=1 m=1

R1 VDD mn {latch1_vsw/latch1_iss} m=1
R2 VDD mp {latch1_vsw/latch1_iss} m=1
R3 VDD oin {latch2_vsw/latch2_iss} m=1
R4 VDD oip {latch2_vsw/latch2_iss} m=1

I1 net2 VSS {latch1_iss}
I2 net6 VSS {latch2_iss}
I3 op VSS {sf_iss}
I4 on VSS {sf_iss}

C1 mp VSS {cwire} m=1
C2 mn VSS {cwire} m=1
C3 oip VSS {cwire} m=1
C4 oin VSS {cwire} m=1

.IC V(mp)={vdd}
.IC V(mn)={vdd-latch1_vsw}
.IC V(oip)={vdd-latch2_vsw}
.IC V(oin)={vdd}
.ends
