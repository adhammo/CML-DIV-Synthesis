.param latch1_winp=$latch1_winp
.param latch1_wclk=$latch1_wclk
.param latch1_wlat=$latch1_wlat
.param latch1_nfinp=$latch1_nfinp
.param latch1_nfclk=$latch1_nfclk
.param latch1_nflat=$latch1_nflat
.param latch1_vsw=$latch1_vsw
.param latch1_iss=$latch1_iss
.param latch2_winp=$latch2_winp
.param latch2_wclk=$latch2_wclk
.param latch2_wlat=$latch2_wlat
.param latch2_nfinp=$latch2_nfinp
.param latch2_nfclk=$latch2_nfclk
.param latch2_nflat=$latch2_nflat
.param latch2_vsw=$latch2_vsw
.param latch2_iss=$latch2_iss
.param sf_w=$sf_w
.param sf_nf=$sf_nf
.param sf_iss=$sf_iss
.param vsw_clk=$vsw_clk
.param cm_clk=$cm_clk
.param cwire=$cwire
.param cload=$cload
.param freq=$freq